library verilog;
use verilog.vl_types.all;
entity square_root_vlg_vec_tst is
end square_root_vlg_vec_tst;
