LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.STD_LOGIC_UNSIGNED;

PACKAGE pacoteBodePunha IS
	TYPE MatrizMUX IS ARRAY(15 downto 0) OF std_logic_vector(4 downto 0);
END;