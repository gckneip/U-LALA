library verilog;
use verilog.vl_types.all;
entity five_bits_sub_adder_vlg_vec_tst is
end five_bits_sub_adder_vlg_vec_tst;
